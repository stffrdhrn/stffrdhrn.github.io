* AC analysis of RC circuit
Vin  2 0 AC SIN(0 0.02 440)
R5  2 1 1K		
C1  1 0 4.7uF		
.tran 0.1m 3m
.plot tran v(2), v(1)
.end
